library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;


entity top_level is
		port(clk, reset_bar, Clock_50: in std_logic
			);
end entity;


architecture behave of top_level is






































end architecture behave;